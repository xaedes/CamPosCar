((lp0
I92
aI190
aI287
aI353
aI417
aI508
aI587
aI548
aI410
aI333
aI202
aI96
aI41
aI36
aI37
a(lp1
I540
aI589
aI577
aI529
aI413
aI365
aI201
aI93
aI31
aI31
aI40
aI95
aI193
aI319
aI435
atp2
.